`timescale 1ns / 1ps


module phy_inout #(
    parameter SIG_TYPE_DIFF   = "FALSE",
    parameter DATA_WIDTH      = 8,
    parameter INIT_VALUE      = 0,
    parameter IDELAY_VALUE    = 0,
    parameter OSERDES_CLK_INV = 0,
    parameter REFCLK_FREQ     = 200.0 // IDELAYCTRL clock input frequency in MHz (200.0-2667.0)
)(
    input                       clk_in,
    input                       clk_div_in,
    input                       ref_clk,//200M
    input                       reset,
//    output                      rst_seq_done,
    input                       tri_t,
    input  [DATA_WIDTH - 1 : 0] data_from_fabric,
    output [DATA_WIDTH - 1 : 0] data_to_fabric,
//    output reg                  data_to_fabric_valid,
    inout                       data_to_and_from_pins_p,
    inout                       data_to_and_from_pins_n,   
    output wire  dq_read_internal
);

wire iob_tri_t;
wire iob_din;
wire iob_dout;
wire iserdes_din;
wire fifo_empty;
wire idelayctrl_rdy;

IDELAYCTRL IDELAYCTRL_inst (
    .RDY(idelayctrl_rdy),
    .REFCLK(ref_clk),
    .RST(reset)
);

generate
if(SIG_TYPE_DIFF == "TRUE") begin: io_pin_diff
    IOBUFDS IOBUFDS_inst (
       .O  (iob_dout               ),     // 1-bit output: Buffer output
       .I  (iob_din                ),     // 1-bit input: Buffer input
       .IO (data_to_and_from_pins_p),     // 1-bit inout: Diff_p inout (connect directly to top-level port)
       .IOB(data_to_and_from_pins_n),     // 1-bit inout: Diff_n inout (connect directly to top-level port)
       .T  (iob_tri_t              )      // 1-bit input: 3-state enable input
    );
end else begin: io_pin_se
    IOBUF IOBUF_inst (
       .O (iob_dout               ),   // 1-bit output: Buffer output
       .I (iob_din                ),   // 1-bit input: Buffer input
       .IO(data_to_and_from_pins_p),   // 1-bit inout: Buffer inout (connect directly to top-level port)
       .T (iob_tri_t              )    // 1-bit input: 3-state enable input
    );
end
endgenerate




IDELAYE2 #(
   .CINVCTRL_SEL("FALSE"),               // Invert CTRL input (TRUE/FALSE)
   .DELAY_SRC("IDATAIN"),                // Delay input (IDATAIN, DATAIN)
   .HIGH_PERFORMANCE_MODE("TRUE"),       // Reduced jitter ("TRUE"), reduced power ("FALSE")
   .IDELAY_TYPE("FIXED"),                // FIXED, VARIABLE, or VAR_LOADABLE
   .IDELAY_VALUE(IDELAY_VALUE),          // Input delay tap setting

   .REFCLK_FREQUENCY(REFCLK_FREQ),       // Reference clock frequency for IDELAYCTRL in MHz (200.0 recommended)
   .SIGNAL_PATTERN("DATA")               // "DATA" for normal signals, "CLOCK" for clock signals
)
IDELAYE2_inst (
   .CNTVALUEOUT(),         // 5-bit output: Counter value output
   .DATAOUT    (iserdes_din), // 1-bit output: Delayed data output
   .C          (clk_div_in),  // 1-bit input: Clock input
   .CE         (1'b0),         // 1-bit input: Enable increment/decrement
   .CINVCTRL   (1'b0),         // 1-bit input: Dynamic clock inversion
   .CNTVALUEIN (5'h0),         // 5-bit input: Counter value input
   .DATAIN     (1'b0),         // 1-bit input: Data input (bypassed in IDATAIN mode)
   .IDATAIN    (iob_dout),     // 1-bit input: Data input from IOB
   .INC        (1'b0),         // 1-bit input: Increment / Decrement tap delay
   .LD         (1'b0),         // 1-bit input: Load IDELAY_VALUE
   .LDPIPEEN   (1'b0),         // 1-bit input: Enable pipeline delay
   .REGRST     (1'b0)          // 1-bit input: Asynchronous Reset
);




ISERDESE2 #(
    .DATA_RATE("DDR"),                   // DDR ģʽ
    .DATA_WIDTH(DATA_WIDTH),             // �������ݿ�� (4 �� 8)
    .INTERFACE_TYPE("NETWORKING"),       // ����Ϊ NETWORKING ģʽ
    .NUM_CE(1),                          // ʹ��һ��ʱ��ʹ��
    .SERDES_MODE("MASTER"),              // ��ģʽ
    .INIT_Q1(1'b0),                      // Q1 �ĳ�ʼֵ
    .INIT_Q2(1'b0),                      // Q2 �ĳ�ʼֵ
    .INIT_Q3(1'b0),                      // Q3 �ĳ�ʼֵ
    .INIT_Q4(1'b0),                      // Q4 �ĳ�ʼֵ
    .SRVAL_Q1(1'b0),                     // ��λֵ
    .SRVAL_Q2(1'b0),
    .SRVAL_Q3(1'b0),
    .SRVAL_Q4(1'b0)
) ISERDESE2_inst (
    .Q1(data_to_fabric[7]),              // �����������λ 1
    .Q2(data_to_fabric[6]),              // �����������λ 2
    .Q3(data_to_fabric[5]),              // �����������λ 3
    .Q4(data_to_fabric[4]),              // �����������λ 4
    .Q5(data_to_fabric[3]),              // �����������λ 5
    .Q6(data_to_fabric[2]),              // �����������λ 6
    .Q7(data_to_fabric[1]),              // �����������λ 7
    .Q8(data_to_fabric[0]),              // �����������λ 8
    .BITSLIP(1'b0),                      // Bit-slip ʹ��
    .CE1(1'b1),                          // ʱ��ʹ��
    .CE2(1'b0),                          // ��ʹ�õڶ�ʹ��
    .CLK(clk_in),                        // ����ʱ������
    .CLKB(~clk_in),                      // �������ʱ�� (UltraScale �� `CLK_B`)
    .CLKDIV(clk_div_in),                 // ��Ƶ���ʱ��
    .DDLY(1'b0), // ? �ӳٺ���ź��� DDLY
    .D(iob_dout),            // D �ڿ��ţ���0
    .RST(reset),                         // �첽��λ
    .SHIFTIN1(1'b0),                     // �������� (δʹ��)
    .SHIFTIN2(1'b0),                     // �������� (δʹ��)
    .SHIFTOUT1(),                        // ������� (δʹ��)
    .SHIFTOUT2()                         // ������� (δʹ��)
);

// OSERDESE2: ���������ģ��
// ����: ������FPGA�ڲ��߼��Ĳ�������(data_from_fabric)ת���ɸ��ٴ���������(iob_din)����ͨ��IO���ŷ��ͳ�ȥ��
//       ͬʱ����Ҳ����IO���ŵ���̬ʹ���ź�(iob_tri_t)��
OSERDESE2 #(
    // --- �������� ---
    .DATA_RATE_OQ("DDR"),      // �������(OQ)ʹ��˫����������(DDR)����CLK�������غ��½��ض���������
    .DATA_RATE_TQ("SDR"),      // ��̬����(TQ)ʹ�õ�����������(SDR)����CLKDIV�������ر仯��ȷ���ź��ȶ�
    .DATA_WIDTH(8),            // �������������λ��Ϊ8λ (D1-D8)
    .INIT_OQ(1'b0),            // OQ�˿ڳ�ʼֵΪ0
    .INIT_TQ(1'b0),            // TQ�˿ڳ�ʼֵΪ0
    .SERDES_MODE("MASTER"),    // ����ΪMASTERģʽ����Ϊ�����Ĵ�����ʹ��
    .SRVAL_OQ(1'b0),           // ��λʱOQ�˿ڵ�ֵ
    .SRVAL_TQ(1'b0),           // ��λʱTQ�˿ڵ�ֵ
    .TRISTATE_WIDTH(1)         // ��̬�����źŵĿ��
) OSERDESE2_inst (
    // --- ����˿� ---
    .OQ    (iob_din),          // ����������������ӵ�IOBUF�������
    .TQ    (iob_tri_t),        // ��̬�����ź���������ӵ�IOBUF����̬ʹ�ܶ�
    // --- ʱ�Ӻ͸�λ ---
    .CLK   (clk_in),           // ���ٴ���ʱ��
    .CLKDIV(clk_div_in),       // ���ٲ���ʱ�� (����FPGA�߼�)
    .RST   (reset),            // �첽��λ�ź�
    // --- ������������ ---
    .D1    (data_from_fabric[0]), // ������������λ1
    .D2    (data_from_fabric[1]),
    .D3    (data_from_fabric[2]),
    .D4    (data_from_fabric[3]),
    .D5    (data_from_fabric[4]),
    .D6    (data_from_fabric[5]),
    .D7    (data_from_fabric[6]),
    .D8    (data_from_fabric[7]),
    .OCE   (1'b1),             // ���ʱ��ʹ�ܣ��ߵ�ƽ��Ч
    // --- ��̬�������� ---
    .T1    (tri_t),            // ��̬���������źţ������ϲ��߼�
    .T2    (),                 // δʹ�õ���̬��������
    .T3    (),
    .T4    (),
    .TCE   (1'b1),             // ��̬����ʱ��ʹ�ܣ��ߵ�ƽ��Ч
    // --- �����˿� (δʹ��) ---
    .SHIFTIN1(1'b0),
    .SHIFTIN2(1'b0),
    .SHIFTOUT1(),
    .SHIFTOUT2()
);

assign dq_read_internal = iob_dout;
assign dq_read_interna2 = ~dq_read_internal;

endmodule
